//用于根据指令的op部分和func部分产生对应的内部控制信号
module cpu_control_single(
    input [5:0] op,//每条指令开头的6位op部分
    input [5:0] fun,//R类型的fun部分
    input z,//zero
    output wmem,//写内存使能
    output wreg,//写寄存器使能
    output regrt,
    output m2reg,//从内存读数据到寄存器
    output [3:0]aluc,//alu的选择码
    output shift,//移位
    output aluimm,//立即数
    output [1:0]pcsource,//下一个PC的选择码
    output jal_c,
    output sext
);

wire type = ~|op;
wire add_c = type & fun[5] & ~fun[4] & ~fun[3] & ~fun[2] & ~fun[1] & ~fun[0];
wire sub_c = type & fun[5] & ~fun[4] & ~fun[3] & ~fun[2] & fun[1] & ~fun[0];
wire and_c = type & fun[5] & ~fun[4] & ~fun[3] & fun[2] & ~fun[1] & ~fun[0];
wire or_c =  type & fun[5] & ~fun[4] & ~fun[3] & fun[2] & ~fun[1] & fun[0];
wire xor_c = type & fun[5] & ~fun[4] & ~fun[3] & fun[2] & fun[1] & ~fun[0];
wire sll_c = type & ~fun[5] & ~fun[4] & ~fun[3] & ~fun[2] & ~fun[1] & ~fun[0];
wire srl_c = type & ~fun[5] & ~fun[4] & ~fun[3] & ~fun[2] & fun[1] & ~fun[0];
wire sra_c =  type & ~fun[5] & ~fun[4] & ~fun[3] & ~fun[2] & fun[1] & fun[0];
wire jr_c = type & ~fun[5] & ~fun[4] & fun[3] & ~fun[2] & ~fun[1] & ~fun[0];

wire addi = ~op[5] & ~op[4] & op[3] & ~op[2] & ~op[1] & ~op[0];
wire andi = ~op[5] & ~op[4] & op[3] & op[2] & ~op[1] & ~op[0];
wire ori = ~op[5] & ~op[4] & op[3] & op[2] & ~op[1] & op[0];
wire xori = ~op[5] & ~op[4] & op[3] & op[2] & op[1] & ~op[0];

wire lw_c = op[5] & ~op[4] & ~op[3] & ~op[2] & op[1] & op[0];
wire sw_c = op[5] & ~op[4] & op[3] & ~op[2] & op[1] & op[0];

wire beq_c = ~op[5] & ~op[4] & ~op[3] & op[2] & ~op[1] & ~op[0];
wire bne_c = ~op[5] & ~op[4] & ~op[3] & op[2] & ~op[1] & op[0];
wire lui_c = ~op[5] & ~op[4] & op[3] & op[2] & op[1] & op[0];
wire j_c = ~op[5] & ~op[4] & ~op[3] & ~op[2] & op[1] & ~op[0];


assign jal_c = ~op[5] & ~op[4] & ~op[3] & ~op[2] & op[1] & op[0];
assign wreg = add_c | sub_c | and_c | or_c | xor_c | sll_c | srl_c | sra_c | addi | andi | ori | xori | lw_c | lui_c | jal_c;
assign regrt = addi | andi | ori | xori | lw_c | lui_c | jal_c; 
assign m2reg = lw_c;
assign shift = sll_c | srl_c | sra_c;
assign aluimm = addi | andi | ori | xori |lw_c | lui_c | sw_c;
assign sext = addi | lw_c | sw_c | beq_c | bne_c;
assign aluc = {sra_c,{sub_c | or_c | srl_c | sra_c | ori | lui_c},{xor_c | sll_c | srl_c | sra_c | xori | beq_c | bne_c | lui_c},{and_c | or_c | sll_c | srl_c | sra_c | andi | ori}};
assign wmem = sw_c;
assign pcsource[1] = jr_c | j_c | jal_c;
assign pcsource[0] = (beq_c & z) | (bne_c & ~z) | j_c | jal_c;
//assign pcsource = {{jr_c | j_c | jal_c},{beq_c & z | bne_c & ~z | j_c | jal_c}};

endmodule 